$readmemh("new_code0.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[0].RAM.Mem);
$readmemh("new_code1.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[1].RAM.Mem);
$readmemh("new_code2.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[2].RAM.Mem);
$readmemh("new_code3.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[3].RAM.Mem);
$readmemh("new_code4.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[4].RAM.Mem);
$readmemh("new_code5.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[5].RAM.Mem);
$readmemh("new_code6.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[6].RAM.Mem);
$readmemh("new_code7.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[7].RAM.Mem);
$readmemh("new_code8.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[8].RAM.Mem);
$readmemh("new_code9.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[9].RAM.Mem);
$readmemh("new_code10.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[10].RAM.Mem);
$readmemh("new_code11.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[11].RAM.Mem);
$readmemh("new_code12.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[12].RAM.Mem);
$readmemh("new_code13.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[13].RAM.Mem);
$readmemh("new_code14.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[14].RAM.Mem);
$readmemh("new_code15.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[15].RAM.Mem);
$readmemh("new_code16.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[16].RAM.Mem);
$readmemh("new_code17.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[17].RAM.Mem);
$readmemh("new_code18.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[18].RAM.Mem);
$readmemh("new_code19.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[19].RAM.Mem);
$readmemh("new_code20.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[20].RAM.Mem);
$readmemh("new_code21.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[21].RAM.Mem);
$readmemh("new_code22.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[22].RAM.Mem);
$readmemh("new_code23.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[23].RAM.Mem);
$readmemh("new_code24.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[24].RAM.Mem);
$readmemh("new_code25.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[25].RAM.Mem);
$readmemh("new_code26.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[26].RAM.Mem);
$readmemh("new_code27.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[27].RAM.Mem);
$readmemh("new_code28.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[28].RAM.Mem);
$readmemh("new_code29.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[29].RAM.Mem);
$readmemh("new_code30.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[30].RAM.Mem);
$readmemh("new_code31.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[31].RAM.Mem);
$readmemh("new_code32.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[32].RAM.Mem);
$readmemh("new_code33.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[33].RAM.Mem);
$readmemh("new_code34.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[34].RAM.Mem);
$readmemh("new_code35.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[35].RAM.Mem);
$readmemh("new_code36.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[36].RAM.Mem);
$readmemh("new_code37.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[37].RAM.Mem);
$readmemh("new_code38.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[38].RAM.Mem);
$readmemh("new_code39.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[39].RAM.Mem);
$readmemh("new_code40.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[40].RAM.Mem);
$readmemh("new_code41.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[41].RAM.Mem);
$readmemh("new_code42.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[42].RAM.Mem);
$readmemh("new_code43.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[43].RAM.Mem);
$readmemh("new_code44.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[44].RAM.Mem);
$readmemh("new_code45.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[45].RAM.Mem);
$readmemh("new_code46.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[46].RAM.Mem);
$readmemh("new_code47.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[47].RAM.Mem);
$readmemh("new_code48.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[48].RAM.Mem);
$readmemh("new_code49.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[49].RAM.Mem);
$readmemh("new_code50.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[50].RAM.Mem);
$readmemh("new_code51.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[51].RAM.Mem);
$readmemh("new_code52.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[52].RAM.Mem);
$readmemh("new_code53.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[53].RAM.Mem);
$readmemh("new_code54.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[54].RAM.Mem);
$readmemh("new_code55.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[55].RAM.Mem);
$readmemh("new_code56.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[56].RAM.Mem);
$readmemh("new_code57.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[57].RAM.Mem);
$readmemh("new_code58.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[58].RAM.Mem);
$readmemh("new_code59.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[59].RAM.Mem);
$readmemh("new_code60.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[60].RAM.Mem);
$readmemh("new_code61.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[61].RAM.Mem);
$readmemh("new_code62.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[62].RAM.Mem);
$readmemh("new_code63.mem", mb_wrapper_tb.mb_wrapper.mb_i.axi_oram_0.inst.fake_mig.synth_dram.RAM_BLOCK[63].RAM.Mem);
