
//==============================================================================
//	Section:	Includes
//==============================================================================
`include "Const.vh"
//==============================================================================

`timescale 1ns/1ns

//==============================================================================
//	Module:		testUARTTop
//	Desc:		Works for VC707 & KC705
//==============================================================================
module testUARTTop(
			output	[7:0]	led,

			input			sys_clk_p,
			input			sys_clk_n,
			input			sys_rst,

			output			uart_txd,
			input			uart_rxd
	);
	
	//------------------------------------------------------------------------------
	//	Wires & Regs
	//------------------------------------------------------------------------------

    wire  					Clock_Bufg, Clock;
	
	//------------------------------------------------------------------------------
	//	Clocking
	//------------------------------------------------------------------------------
		
    IBUFGDS		ibufgds(	.I(						sys_clk_p),
							.IB(					sys_clk_n),
							.O(						Clock_Bufg));
    BUFG		bufg(		.I(						Clock_Bufg),
							.O(						Clock));
		
	//------------------------------------------------------------------------------
	// 	Loopback test
	//------------------------------------------------------------------------------
	
	UARTLoopback	cut(	.Clock(					Clock), 
							.Reset(					sys_rst),
							.UARTTX(				uart_txd),	
							.UARTRX(				uart_rxd),
							.LastWord(				led));
	
	//------------------------------------------------------------------------------
endmodule
//------------------------------------------------------------------------------